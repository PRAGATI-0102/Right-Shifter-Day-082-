`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 07/01/2023 12:19:32 AM
// Design Name: 
// Module Name: right_shift
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module right_shift(
      input clk, rst,
	  input [3:0] din,
	  output reg [3:0] dout);

	always @(posedge clk or posedge rst) 
	begin
	  if (rst) 
          begin
            dout <= 4'b0000;
          end
	  else 
          begin
            dout[0] <= din[0];
            dout <= {1'b0, din[3:1]};    
          end
	end
endmodule
